

module multiple_echo (sysclk, data_in, data_out, data_valid);

	input				sysclk;		// system clock
	input [9:0]		data_in;		// 10-bit input data
	input 			data_valid;	// asserted when sample data is ready for processing
	output [9:0] 	data_out;	// 10-bit output data

	wire				sysclk ;
	wire [9:0]		data_in;
	reg [9:0] 		data_out;
	wire [9:0]		x,q,y;
	wire full; 
	
	parameter 		ADC_OFFSET = 10'd512;
	parameter 		DAC_OFFSET = 10'd512;

	assign x = data_in[9:0] - ADC_OFFSET;		// x is input in 2's complement
	
	// This part should include your own processing hardware 
	// ... that takes x to produce y
	// ... In this case, it is ALL PASS.
 
	pulse_gen  PULSE (wren, data_valid, sysclk); 
	fifo_fsm fsm(sysclk, full, fifo_state); 
	FIFO fifo(sysclk, y, fifo_state&&wren, wren,full, q);
	assign y = x - {q[9],q[9:1]}; 
	
	//  Now clock y output with system clock
	always @(posedge sysclk)
		if (wren == 1'b1)
			data_out <= y + DAC_OFFSET;  
		 
endmodule
	